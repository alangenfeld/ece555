`timescale 1ns / 1ns 
module cds_alias(output o, input i );
assign o =i;

endmodule
