module fsm(input clk, rst,
    output reg [4:0] rd_enA, rd_enB, wr_en,
    output reg done, ERROR);


   



endmodule; // fsm
