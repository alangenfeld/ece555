// Library - ece555_final, Cell - Shifter_4_32, View - schematic
// LAST TIME SAVED: Dec  4 17:01:22 2010
// NETLIST TIME: Dec  7 19:22:19 2010
`timescale 1ns / 1ns 

module Shifter_4_32 ( OUT, IN, LEFT_NOT, L_SHIFT, NO_SHIFT, OLD_NOT,
     RIGHT_NOT, R_SHIFT );

input  LEFT_NOT, L_SHIFT, NO_SHIFT, OLD_NOT, RIGHT_NOT, R_SHIFT;

output [31:0]  OUT;

input [31:0]  IN;


specify 
    specparam CDS_LIBNAME  = "ece555_final";
    specparam CDS_CELLNAME = "Shifter_4_32";
    specparam CDS_VIEWNAME = "schematic";
endspecify

lr_1b I260 ( OUT[31], IN[27], L_SHIFT, NO_SHIFT, IN[31],
     0, R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I259 ( OUT[30], IN[26], L_SHIFT, NO_SHIFT, IN[30],
     0, R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I258 ( OUT[29], IN[25], L_SHIFT, NO_SHIFT, IN[29],
     0, R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I257 ( OUT[28], IN[24], L_SHIFT, NO_SHIFT, IN[28],
     0, R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I256 ( OUT[24], IN[20], L_SHIFT, NO_SHIFT, IN[24], IN[28],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I255 ( OUT[25], IN[21], L_SHIFT, NO_SHIFT, IN[25], IN[29],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I254 ( OUT[26], IN[22], L_SHIFT, NO_SHIFT, IN[26], IN[30],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I253 ( OUT[27], IN[23], L_SHIFT, NO_SHIFT, IN[27], IN[31],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I252 ( OUT[19], IN[15], L_SHIFT, NO_SHIFT, IN[19], IN[23],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I251 ( OUT[18], IN[14], L_SHIFT, NO_SHIFT, IN[18], IN[22],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I250 ( OUT[17], IN[13], L_SHIFT, NO_SHIFT, IN[17], IN[21],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I249 ( OUT[16], IN[12], L_SHIFT, NO_SHIFT, IN[16], IN[20],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I248 ( OUT[20], IN[16], L_SHIFT, NO_SHIFT, IN[20], IN[24],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I247 ( OUT[21], IN[17], L_SHIFT, NO_SHIFT, IN[21], IN[25],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I246 ( OUT[22], IN[18], L_SHIFT, NO_SHIFT, IN[22], IN[26],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I245 ( OUT[23], IN[19], L_SHIFT, NO_SHIFT, IN[23], IN[27],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I244 ( OUT[7], IN[3], L_SHIFT, NO_SHIFT, IN[7], IN[11], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I243 ( OUT[6], IN[2], L_SHIFT, NO_SHIFT, IN[6], IN[10], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I242 ( OUT[5], IN[1], L_SHIFT, NO_SHIFT, IN[5], IN[9], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I241 ( OUT[4], IN[0], L_SHIFT, NO_SHIFT, IN[4], IN[8], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I240 ( OUT[0], 0, L_SHIFT, NO_SHIFT, IN[0], IN[4],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I239 ( OUT[1], 0, L_SHIFT, NO_SHIFT, IN[1], IN[5],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I238 ( OUT[2], 0, L_SHIFT, NO_SHIFT, IN[2], IN[6],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I237 ( OUT[3], 0, L_SHIFT, NO_SHIFT, IN[3], IN[7],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I236 ( OUT[8], IN[4], L_SHIFT, NO_SHIFT, IN[8], IN[12], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I235 ( OUT[9], IN[5], L_SHIFT, NO_SHIFT, IN[9], IN[13], R_SHIFT,
     LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I234 ( OUT[10], IN[6], L_SHIFT, NO_SHIFT, IN[10], IN[14],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I233 ( OUT[11], IN[7], L_SHIFT, NO_SHIFT, IN[11], IN[15],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I232 ( OUT[12], IN[8], L_SHIFT, NO_SHIFT, IN[12], IN[16],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I231 ( OUT[13], IN[9], L_SHIFT, NO_SHIFT, IN[13], IN[17],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I230 ( OUT[14], IN[10], L_SHIFT, NO_SHIFT, IN[14], IN[18],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);
lr_1b I229 ( OUT[15], IN[11], L_SHIFT, NO_SHIFT, IN[15], IN[19],
     R_SHIFT, LEFT_NOT, OLD_NOT, RIGHT_NOT);

endmodule
